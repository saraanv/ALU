library verilog;
use verilog.vl_types.all;
entity prj_vlg_vec_tst is
end prj_vlg_vec_tst;
